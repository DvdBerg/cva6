/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the "License"); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [63:0]  addr_i,
   output logic [63:0]  rdata_o
);
    localparam int RomSize = 855;

    const logic [RomSize-1:0][63:0] mem = {
        64'h00000000_00000000,
        64'h0a0d2165_6e6f6420,
        64'h00000000_00206567,
        64'h616d6920_746f6f62,
        64'h20676e69_79706f63,
        64'h00000000_00000009,
        64'h3a656d61_6e090a0d,
        64'h00093a73_65747562,
        64'h69727474_61090a0d,
        64'h00000009_3a61626c,
        64'h20747361_6c090a0d,
        64'h0000093a_61626c20,
        64'h74737269_66090a0d,
        64'h00000000_00000000,
        64'h09202020_20203a64,
        64'h69756720_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_00000000,
        64'h093a6469_75672065,
        64'h70797420_6e6f6974,
        64'h69747261_70090a0d,
        64'h00000000_20797274,
        64'h6e65206e_6f697469,
        64'h74726170_20747067,
        64'h00000009_20203a73,
        64'h65697274_6e65206e,
        64'h6f697469_74726170,
        64'h20657a69_73090a0d,
        64'h00000009_3a736569,
        64'h72746e65_206e6f69,
        64'h74697472_61702072,
        64'h65626d75_6e090a0d,
        64'h00000009_2020203a,
        64'h61626c20_73656972,
        64'h746e6520_6e6f6974,
        64'h69747261_70090a0d,
        64'h00093a61_646c2070,
        64'h756b6361_62090a0d,
        64'h00000000_00000000,
        64'h093a6162_6c20746e,
        64'h65727275_63090a0d,
        64'h00000009_3a646576,
        64'h72657365_72090a0d,
        64'h00093a72_65646165,
        64'h685f6372_63090a0d,
        64'h00000000_00000909,
        64'h3a657a69_73090a0d,
        64'h00000009_3a6e6f69,
        64'h73697665_72090a0d,
        64'h0000093a_65727574,
        64'h616e6769_73090a0d,
        64'h00000000_003a7265,
        64'h64616568_20656c62,
        64'h6174206e_6f697469,
        64'h74726170_20747067,
        64'h0000203a_65756c61,
        64'h76206e72_75746572,
        64'h2079706f_63206473,
        64'h00000000_0000000a,
        64'h0d216465_6c696166,
        64'h20647261_63204453,
        64'h00000000_0000000a,
        64'h0d216465_7a696c61,
        64'h6974696e_69206473,
        64'h00000000_0a0d676e,
        64'h69746978_65202e2e,
        64'h2e647320_657a696c,
        64'h61697469_6e692074,
        64'h6f6e2064_6c756f63,
        64'h00000000_0000002e,
        64'h00000000_0000000a,
        64'h0d6b636f_6c622044,
        64'h53206461_65722074,
        64'h6f6e2064_6c756f63,
        64'h0000000a_0d202e2e,
        64'h2e445320_676e697a,
        64'h696c6169_74696e69,
        64'h00000031_34646d63,
        64'h00000035_35646d63,
        64'h00000000_30646d63,
        64'h00000020_3a206573,
        64'h6e6f7073_65720920,
        64'h00000000_0020646e,
        64'h616d6d6f_63204453,
        64'h00000000_203f3f79,
        64'h74706d65_20746f6e,
        64'h206f6669_66207872,
        64'h00000000_00000a0d,
        64'h2164657a_696c6169,
        64'h74696e69_20495053,
        64'h00000000_00007830,
        64'h203a7375_74617473,
        64'h00000000_00000a0d,
        64'h49505320_74696e69,
        64'h00000a0d_21646c72,
        64'h6f57206f_6c6c6548,
        64'h00322d74_6c756166,
        64'h65642d69_72742c78,
        64'h6e6c7800_746c7561,
        64'h6665642d_6972742c,
        64'h786e6c78_006c6175,
        64'h642d7369_2c786e6c,
        64'h7800746e_65736572,
        64'h702d7470_75727265,
        64'h746e692c_786e6c78,
        64'h00687464_69772d32,
        64'h6f697067_2c786e6c,
        64'h78006874_6469772d,
        64'h6f697067_2c786e6c,
        64'h7800322d_746c7561,
        64'h6665642d_74756f64,
        64'h2c786e6c_7800746c,
        64'h75616665_642d7475,
        64'h6f642c78_6e6c7800,
        64'h322d7374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007374_75706e69,
        64'h2d6c6c61_2c786e6c,
        64'h78007265_6c6c6f72,
        64'h746e6f63_2d6f6970,
        64'h6700736c_6c65632d,
        64'h6f697067_23007077,
        64'h2d656c62_61736964,
        64'h00736567_6e61722d,
        64'h65676174_6c6f7600,
        64'h79636e65_75716572,
        64'h662d7861_6d2d6970,
        64'h73006f69_7461722d,
        64'h6b63732c_786e6c78,
        64'h00737469_622d7265,
        64'h66736e61_72742d6d,
        64'h756e2c78_6e6c7800,
        64'h73746962_2d73732d,
        64'h6d756e2c_786e6c78,
        64'h00747369_78652d6f,
        64'h6669662c_786e6c78,
        64'h00796c69_6d61662c,
        64'h786e6c78_00687464,
        64'h69772d6f_692d6765,
        64'h72007466_6968732d,
        64'h67657200_73747075,
        64'h72726574_6e690074,
        64'h6e657261_702d7470,
        64'h75727265_746e6900,
        64'h64656570_732d746e,
        64'h65727275_63007665,
        64'h646e2c76_63736972,
        64'h00797469_726f6972,
        64'h702d7861_6d2c7663,
        64'h73697200_73656d61,
        64'h6e2d6765_72006465,
        64'h646e6574_78652d73,
        64'h74707572_7265746e,
        64'h69007365_676e6172,
        64'h00646564_6e657073,
        64'h75732d65_74617473,
        64'h2d6e6961_74657200,
        64'h72656767_6972742d,
        64'h746c7561_6665642c,
        64'h78756e69_6c00736f,
        64'h69706700_656c646e,
        64'h61687000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h00736c6c_65632d74,
        64'h70757272_65746e69,
        64'h23007469_6c70732d,
        64'h626c7400_65707974,
        64'h2d756d6d_00617369,
        64'h2c766373_69720073,
        64'h75746174_73006765,
        64'h72006570_79745f65,
        64'h63697665_64007963,
        64'h6e657571_6572662d,
        64'h6b636f6c_63007963,
        64'h6e657571_6572662d,
        64'h65736162_656d6974,
        64'h00687461_702d7475,
        64'h6f647473_006c6564,
        64'h6f6d0065_6c626974,
        64'h61706d6f_6300736c,
        64'h6c65632d_657a6973,
        64'h2300736c_6c65632d,
        64'h73736572_64646123,
        64'h09000000_02000000,
        64'h02000000_02000000,
        64'h01000000_b5000000,
        64'h04000000_03000000,
        64'hffffffff_ad020000,
        64'h04000000_03000000,
        64'hffffffff_9c020000,
        64'h04000000_03000000,
        64'h01000000_8f020000,
        64'h04000000_03000000,
        64'h00000000_78020000,
        64'h04000000_03000000,
        64'h08000000_67020000,
        64'h04000000_03000000,
        64'h08000000_57020000,
        64'h04000000_03000000,
        64'h00000000_43020000,
        64'h04000000_03000000,
        64'h00000000_31020000,
        64'h04000000_03000000,
        64'h00000000_1f020000,
        64'h04000000_03000000,
        64'h00000000_0f020000,
        64'h04000000_03000000,
        64'h00000100_00000000,
        64'h00000040_00000000,
        64'h67000000_10000000,
        64'h03000000_ff010000,
        64'h00000000_03000000,
        64'h00000000_612e3030,
        64'h2e312d6f_6970672d,
        64'h7370782c_786e6c78,
        64'h1b000000_15000000,
        64'h03000000_02000000,
        64'hf3010000_04000000,
        64'h03000000_00000030,
        64'h30303030_30303440,
        64'h6f697067_01000000,
        64'h02000000_02000000,
        64'he8010000_00000000,
        64'h03000000_e40c0000,
        64'he40c0000_d9010000,
        64'h08000000_03000000,
        64'h20bcbe00_c7010000,
        64'h04000000_03000000,
        64'h00000000_67000000,
        64'h04000000_03000000,
        64'h00000000_746f6c73,
        64'h2d697073_2d636d6d,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h40636d6d_01000000,
        64'h04000000_b8010000,
        64'h04000000_03000000,
        64'h08000000_a1010000,
        64'h04000000_03000000,
        64'h01000000_90010000,
        64'h04000000_03000000,
        64'h01000000_80010000,
        64'h04000000_03000000,
        64'h00377865_746e696b,
        64'h74010000_08000000,
        64'h03000000_00100000,
        64'h00000000_00000020,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h02000000_02000000,
        64'h52010000_08000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00000000,
        64'h0f000000_04000000,
        64'h03000000_01000000,
        64'h00000000_04000000,
        64'h03000000_00612e30,
        64'h302e322d_6970732d,
        64'h7370782c_786e6c78,
        64'h00622e30_302e322d,
        64'h6970732d_7370782c,
        64'h786e6c78_1b000000,
        64'h28000000_03000000,
        64'h00000000_30303030,
        64'h30303032_40697073,
        64'h2d737078_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h03000000_41010000,
        64'h04000000_03000000,
        64'h00100000_00000000,
        64'h00000018_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h06000000_05000000,
        64'h04000000_52010000,
        64'h10000000_03000000,
        64'h00007265_6d69745f,
        64'h6270612c_706c7570,
        64'h1b000000_0f000000,
        64'h03000000_00003030,
        64'h30303030_38314072,
        64'h656d6974_01000000,
        64'h02000000_04000000,
        64'h67010000_04000000,
        64'h03000000_02000000,
        64'h5d010000_04000000,
        64'h03000000_01000000,
        64'h52010000_04000000,
        64'h03000000_03000000,
        64'h41010000_04000000,
        64'h03000000_00c20100,
        64'h33010000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00100000,
        64'h00000000_00000010,
        64'h00000000_67000000,
        64'h10000000_03000000,
        64'h00303537_3631736e,
        64'h1b000000_08000000,
        64'h03000000_00000030,
        64'h30303030_30303140,
        64'h74726175_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00100000_00000000,
        64'h00000000_00000000,
        64'h67000000_10000000,
        64'h03000000_ffff0000,
        64'h02000000_f7000000,
        64'h08000000_03000000,
        64'h00333130_2d677562,
        64'h65642c76_63736972,
        64'h1b000000_10000000,
        64'h03000000_00003040,
        64'h72656c6c_6f72746e,
        64'h6f632d67_75626564,
        64'h01000000_02000000,
        64'h03000000_b5000000,
        64'h04000000_03000000,
        64'h1e000000_28010000,
        64'h04000000_03000000,
        64'h07000000_15010000,
        64'h04000000_03000000,
        64'h00000004_00000000,
        64'h0000000c_00000000,
        64'h67000000_10000000,
        64'h03000000_09000000,
        64'h02000000_0b000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'ha0000000_00000000,
        64'h03000000_00306369,
        64'h6c702c76_63736972,
        64'h1b000000_0c000000,
        64'h03000000_01000000,
        64'h8f000000_04000000,
        64'h03000000_00000000,
        64'h00000000_04000000,
        64'h03000000_00000000,
        64'h30303030_30306340,
        64'h72656c6c_6f72746e,
        64'h6f632d74_70757272,
        64'h65746e69_01000000,
        64'h02000000_006c6f72,
        64'h746e6f63_0b010000,
        64'h08000000_03000000,
        64'h00000c00_00000000,
        64'h00000002_00000000,
        64'h67000000_10000000,
        64'h03000000_07000000,
        64'h02000000_03000000,
        64'h02000000_f7000000,
        64'h10000000_03000000,
        64'h00000000_30746e69,
        64'h6c632c76_63736972,
        64'h1b000000_0d000000,
        64'h03000000_00000030,
        64'h30303030_30324074,
        64'h6e696c63_01000000,
        64'hf0000000_00000000,
        64'h03000000_00007375,
        64'h622d656c_706d6973,
        64'h00636f73_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h1f000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00636f73_01000000,
        64'h02000000_02000000,
        64'hd9000000_00000000,
        64'h03000000_00000074,
        64'h61656274_72616568,
        64'hc3000000_0a000000,
        64'h03000000_00000000,
        64'h01000000_01000000,
        64'hbd000000_0c000000,
        64'h03000000_00000064,
        64'h656c2d74_61656274,
        64'h72616568_01000000,
        64'h00000073_64656c2d,
        64'h6f697067_1b000000,
        64'h0a000000_03000000,
        64'h00000000_7364656c,
        64'h01000000_02000000,
        64'h0000003c_00000000,
        64'h00000080_00000000,
        64'h67000000_10000000,
        64'h03000000_00007972,
        64'h6f6d656d_5b000000,
        64'h07000000_03000000,
        64'h00303030_30303030,
        64'h38407972_6f6d656d,
        64'h01000000_02000000,
        64'h02000000_02000000,
        64'h02000000_b5000000,
        64'h04000000_03000000,
        64'h00006374_6e692d75,
        64'h70632c76_63736972,
        64'h1b000000_0f000000,
        64'h03000000_a0000000,
        64'h00000000_03000000,
        64'h01000000_8f000000,
        64'h04000000_03000000,
        64'h00000000_72656c6c,
        64'h6f72746e_6f632d74,
        64'h70757272_65746e69,
        64'h01000000_85000000,
        64'h00000000_03000000,
        64'h00003933_76732c76,
        64'h63736972_7c000000,
        64'h0b000000_03000000,
        64'h00006364_66616d69,
        64'h34367672_72000000,
        64'h0b000000_03000000,
        64'h00000076_63736972,
        64'h00656e61_69726120,
        64'h2c687465_1b000000,
        64'h12000000_03000000,
        64'h00000000_79616b6f,
        64'h6b000000_05000000,
        64'h03000000_00000000,
        64'h67000000_04000000,
        64'h03000000_00757063,
        64'h5b000000_04000000,
        64'h03000000_80f0fa02,
        64'h4b000000_04000000,
        64'h03000000_00000030,
        64'h40757063_01000000,
        64'h40787d01_38000000,
        64'h04000000_03000000,
        64'h00000000_0f000000,
        64'h04000000_03000000,
        64'h01000000_00000000,
        64'h04000000_03000000,
        64'h00000000_73757063,
        64'h01000000_02000000,
        64'h00000030_30323531,
        64'h313a3030_30303030,
        64'h30314074_7261752f,
        64'h636f732f_2c000000,
        64'h1a000000_03000000,
        64'h00006e65_736f6863,
        64'h01000000_00657261,
        64'h622d656e_61697261,
        64'h2c687465_26000000,
        64'h10000000_03000000,
        64'h00766564_2d657261,
        64'h622d656e_61697261,
        64'h2c687465_1b000000,
        64'h14000000_03000000,
        64'h02000000_0f000000,
        64'h04000000_03000000,
        64'h02000000_00000000,
        64'h04000000_03000000,
        64'h00000000_01000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'hc0080000_c0020000,
        64'h00000000_10000000,
        64'h11000000_28000000,
        64'hf8080000_38000000,
        64'hb80b0000_edfe0dd0,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h46454443_42413938,
        64'h37363534_33323130,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_0000a001,
        64'h84021325_85930000,
        64'h0597047e_0010041b,
        64'he909d05f_f0ef057e,
        64'h65a14505_ec0ff0ef,
        64'hd0850513_00001517,
        64'he88ff0ef_e4060805,
        64'h05132005_85931141,
        64'h02faf537_65f1b38d,
        64'hee4ff0ef_01c50513,
        64'h00001517_bbd9d765,
        64'h05130000_1517f7cf,
        64'hf0ef8526_f00ff0ef,
        64'he7850513_00001517,
        64'hf0cff0ef_e6c50513,
        64'h00001517_bbfdd9e5,
        64'h05130000_1517fa4f,
        64'hf0ef8526_f28ff0ef,
        64'hea050513_00001517,
        64'hf34ff0ef_e9450513,
        64'h00001517_c92984aa,
        64'hc3bff0ef_8556865a,
        64'h020ba583_f50ff0ef,
        64'h07050513_00001517,
        64'hf3849de3_08090913,
        64'h080a0993_f68ff0ef,
        64'h2485df25_05130000,
        64'h1517ff3a_1be383ff,
        64'hf0ef0a05_000a4503,
        64'hf84ff0ef_09450513,
        64'h00001517_813ff0ef,
        64'h01093503_f98ff0ef,
        64'h09850513_00001517,
        64'h827ff0ef_00893503,
        64'hfacff0ef_09c50513,
        64'h00001517_83bff0ef,
        64'hfb898a13_00093503,
        64'hfc4ff0ef_0a450513,
        64'h00001517_ff2a1be3,
        64'h899ff0ef_0a05000a,
        64'h4503f909_8a13fe2f,
        64'hf0ef0a25_05130000,
        64'h1517ff9a_19e38b7f,
        64'hf0ef0a05_0007c503,
        64'h014d07b3_4a01803f,
        64'hf0eff809_8d130a65,
        64'h05130000_15178d7f,
        64'hf0ef0ff4_f51381bf,
        64'hf0ef0a25_05130000,
        64'h15174c11_4cc11005,
        64'h1b630201_09130801,
        64'h099384aa_8b8ad31f,
        64'hf0ef850a_46057101,
        64'h04892583_849ff0ef,
        64'hed050513_00001517,
        64'h897ff0ef_455685bf,
        64'hf0ef0c25_05130000,
        64'h15178a9f_f0ef4546,
        64'h86dff0ef_0b450513,
        64'h00001517_8fbff0ef,
        64'h652687ff_f0ef0a65,
        64'h05130000_151790df,
        64'hf0ef7502_891ff0ef,
        64'h0a850513_00001517,
        64'h91fff0ef_65628a3f,
        64'hf0ef0a25_05130000,
        64'h15178f1f_f0ef4552,
        64'h8b5ff0ef_0a450513,
        64'h00001517_903ff0ef,
        64'h45428c7f_f0ef0a65,
        64'h05130000_1517915f,
        64'hf0ef4532_8d9ff0ef,
        64'h0a850513_00001517,
        64'h927ff0ef_45228ebf,
        64'hf0ef0aa5_05130000,
        64'h1517979f_f0ef6502,
        64'h8fdff0ef_0ac50513,
        64'h00001517_909ff0ef,
        64'h09850513_00001517,
        64'hbf5154f9_919ff0ef,
        64'hfa050513_00001517,
        64'h9a7ff0ef_852692bf,
        64'hf0ef0a25_05130000,
        64'h1517937f_f0ef0965,
        64'h05130000_1517c905,
        64'h84aa890a_e3fff0ef,
        64'h850a4585_46057101,
        64'h955ff0ef_09c50513,
        64'h00001517_80826125,
        64'h6d026ca2_6c426be2,
        64'h7b027aa2_7a4279e2,
        64'h690664a6_64468526,
        64'h60e6fa04_011354fd,
        64'h985ff0ef_0a450513,
        64'h00001517_c90ddf1f,
        64'hf0ef8b2e_8aaa1080,
        64'he06ae466_e862ec5e,
        64'hf852fc4e_e0cae4a6,
        64'hec86f05a_f456e8a2,
        64'h711db765_54798082,
        64'h61696baa_6b4a6aea,
        64'h7a0a79aa_794a74ea,
        64'h640e8522_60ae547d,
        64'h9d5ff0ef_0cc50513,
        64'h00001517_c5fff0ef,
        64'hc63ff0ef_c67ff0ef,
        64'hc6bff0ef_c6fff0ef,
        64'hc73ff0ef_c77ff0ef,
        64'hc7bff0ef_a805c81f,
        64'hf0efc8bf_f0ef4531,
        64'h45814605_4401f930,
        64'h45e32004_849319fd,
        64'ha1dff0ef_13450513,
        64'h00001517_e7990359,
        64'he7b30724_1c632901,
        64'h90411442_8c49cb9f,
        64'hf0ef9041_14420085,
        64'h141bcc5f_f0effc94,
        64'h18e30404_0413ff7b,
        64'h15e3892a_f19ff0ef,
        64'h0ff5f593_0b05854a,
        64'h0007c583_016407b3,
        64'h04000b93_4b01c6df,
        64'hf0ef850a_04000593,
        64'h86224901_ff451ee3,
        64'hd03ff0ef_e0048413,
        64'h3e800a93_0fe00a13,
        64'he9592004_8493d1ff,
        64'hf0ef4549_85a20ff6,
        64'h76130016_66130015,
        64'h1613f51f_f0ef0ff4,
        64'h7593f59f_f0ef0ff5,
        64'hf5930084_559bf65f,
        64'hf0ef0ff5_f5930104,
        64'h559bf71f_f0ef4501,
        64'h0184559b_fee79be3,
        64'h078500c6_802300f1,
        64'h06b30800_0713567d,
        64'h47810209_d993842e,
        64'h84aae55e_e95aed56,
        64'hf152f94a_e586fd26,
        64'he1a20206_1993f54e,
        64'h71558082_91411542,
        64'h8d2d8d7d_0055151b,
        64'h17816789_0105551b,
        64'h0105951b_8da900c5,
        64'h95138da9_893d0045,
        64'hd51b8da9_91411542,
        64'h8d5d0522_0085579b,
        64'h808207f5_75138d2d,
        64'h00451593_8d2d0ff5,
        64'h75138d3d_0045d51b,
        64'h0075d79b_8de98082,
        64'h0141853e_640260a2,
        64'h57f5e111_4781f89f,
        64'hf0efc511_57f9efbf,
        64'hf0efc911_57fdeb7f,
        64'hf0effc6d_e07ff0ef,
        64'h347d4429_b91ff0ef,
        64'h27050513_00001517,
        64'hc8bff0ef_e022e406,
        64'h11418082_61050015,
        64'h351364a2_64420004,
        64'h051b60e2_fc940ce3,
        64'he3bff0ef_eb3ff0ef,
        64'h29850513_00001517,
        64'h85aa842a_e55ff0ef,
        64'h02900513_400005b7,
        64'h07700613_fbdff0ef,
        64'h4485e822_ec06e426,
        64'h11018082_01410015,
        64'h3513157d_64020004,
        64'h051b60a2_ef3ff0ef,
        64'h2d250513_85a20000,
        64'h1517e8df_f0ef842a,
        64'he99ff0ef_e022e406,
        64'h03700513_45810650,
        64'h06131141_80826105,
        64'h690264a2_644260e2,
        64'h00153513_f5650513,
        64'h0004051b_01249863,
        64'h88bd00f9_1b634501,
        64'h4785ecdf_f0efed1f,
        64'hf0ef842a_ed7ff0ef,
        64'h84aaeddf_f0efee1f,
        64'hf0efee5f_f0ef892a,
        64'hef1ff0ef_e04ae426,
        64'he822ec06_45211aa0,
        64'h05930870_06131101,
        64'hbfcd4501_80826105,
        64'h690264a2_644260e2,
        64'h4505f89f_f0ef4585,
        64'h36050513_00001517,
        64'hff2495e3_c00df29f,
        64'hf0ef84aa_347df37f,
        64'hf0ef4501_45810950,
        64'h06134905_71040413,
        64'he426ec06_e04a6409,
        64'he8221101_b1f96105,
        64'h35850513_00001517,
        64'h64a260e2_6442da7f,
        64'hf0ef8522_ce9ff0ef,
        64'h3a050513_00001517,
        64'hcf5ff0ef_8526cfbf,
        64'hf0ef842e_e822ec06,
        64'h3a850513_00001517,
        64'h84aae426_11018082,
        64'h61056902_64a26442,
        64'h60e2f47d_147d0007,
        64'hd4634187_d79b0185,
        64'h179bfadf_f0ef0640,
        64'h0413ebbf_f0ef8526,
        64'hec1ff0ef_0ff47513,
        64'hec9ff0ef_0ff57513,
        64'h0084551b_ed5ff0ef,
        64'h0ff57513_0104551b,
        64'hee1ff0ef_0184551b,
        64'hee9ff0ef_04096513,
        64'hfebff0ef_892ae04a,
        64'h84b2842e_e426e822,
        64'hec061101_b7090ff0,
        64'h05138082_557db7d9,
        64'h00d70023_078500f6,
        64'h073306c8_2683ff69,
        64'h8b055178_b77dd6b8,
        64'h07850007_470300f5,
        64'h07338082_4501d3b8,
        64'h4719dbb8_577d2000,
        64'h07b702b6_e1630007,
        64'h869b2000_08372000,
        64'h0537fff5_8b85537c,
        64'h20000737_d3b82000,
        64'h07b71060_0713fff5,
        64'h37fd0001_03200793,
        64'h04b76163_0007871b,
        64'h47812000_06b7dbb8,
        64'h57792000_07b706b7,
        64'hee631000_07938082,
        64'h610564a2_d3b84719,
        64'hdbb86442_0ff47513,
        64'h577d2000_07b760e2,
        64'he25ff0ef_4ac50513,
        64'h00001517_eb3ff0ef,
        64'h91011502_4088e3bf,
        64'hf0ef4ca5_05130000,
        64'h1517e395_8b852401,
        64'h53fc57e0_ff658b05,
        64'h06478493_53f8d3b8,
        64'h10600713_200007b7,
        64'hfff537fd_00010640,
        64'h0793d7a8_dbb85779,
        64'he426e822_ec062000,
        64'h07b71101_bdbd6105,
        64'h4f850513_00001517,
        64'h64a260e2_6442d03c,
        64'h4799e97f_f0ef51e5,
        64'h05130000_1517f25f,
        64'hf0ef9101_02049513,
        64'h2481eaff_f0ef5165,
        64'h05130000_15175064,
        64'hd03c1660_0793ec3f,
        64'hf0ef54a5_05130000,
        64'h1517f51f_f0ef9101,
        64'h02049513_2481edbf,
        64'hf0ef5425_05130000,
        64'h15175064_d03c1040,
        64'h07932000_0437fff5,
        64'h37fd0001_47a9c3b8,
        64'h47292000_07b7f03f,
        64'hf0efe426_e822ec06,
        64'h56250513_11010000,
        64'h15178082_25014108,
        64'h8082c10c_80826105,
        64'h60e2ecff_f0ef0091,
        64'h4503ed7f_f0ef0081,
        64'h4503f55f_f0efec06,
        64'h002c1101_80826145,
        64'h694264e2_740270a2,
        64'hff2410e3_ef9ff0ef,
        64'h00914503_f01ff0ef,
        64'h34610081_4503f81f,
        64'hf0ef0ff5_7513002c,
        64'h0084d533_59610380,
        64'h041384aa_f406e84a,
        64'hec26f022_71798082,
        64'h61456942_64e27402,
        64'h70a2ff24_10e3f3bf,
        64'hf0ef0091_4503f43f,
        64'hf0ef3461_00814503,
        64'hfc3ff0ef_0ff57513,
        64'h002c0084_d53b5961,
        64'h446184aa_f406e84a,
        64'hec26f022_71798082,
        64'h00f58023_0007c783,
        64'h00e580a3_97aa8111,
        64'h00074703_973e00f5,
        64'h771396a7_87930000,
        64'h1797b7f5_0405f93f,
        64'hf0ef8082_01416402,
        64'h60a2e509_00044503,
        64'h842ae406_e0221141,
        64'h808200e7_88230200,
        64'h071300e7_8423fc70,
        64'h071300e7_8623470d,
        64'h00a78223_0ff57513,
        64'h00e78023_0085551b,
        64'h0ff57713_00e78623,
        64'hf8000713_00078223,
        64'h100007b7_02b5553b,
        64'h0045959b_808200a7,
        64'h0023dfe5_0207f793,
        64'h01474783_10000737,
        64'h80820205_75130147,
        64'hc5031000_07b78082,
        64'h0ff57513_00054503,
        64'h808200b5_00238082,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00000000_00000000,
        64'h00048067_01f49493,
        64'h0010049b_b8458593,
        64'h00001597_f1402573,
        64'hff24c6e3_4009091b,
        64'h02000937_00448493,
        64'hfe091ee3_0004a903,
        64'h00092023_00990933,
        64'h00291913_f1402973,
        64'h020004b7_fe090ae3,
        64'h00897913_34402973,
        64'h10500073_ff24c6e3,
        64'h4009091b_02000937,
        64'h00448493_0124a023,
        64'h00100913_020004b7,
        64'h27f000ef_01a11113,
        64'h0210011b_03249663,
        64'hf1402973_00000493,
        64'h30491073_00800913
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    // this prevents spurious Xes from propagating into
    // the speculative fetch stage of the core
    assign rdata_o = (addr_q < RomSize) ? mem[addr_q] : '0;
endmodule
